LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
ENTITY FREQUENCIES IS
	PORT(CLK:IN STD_LOGIC;
		 clk_1k:OUT STD_LOGIC;
		 clk_100hz:out std_logic);
END FREQUENCIES;
ARCHITECTURE BEHAV OF FREQUENCIES IS
BEGIN
	PROCESS(CLK)
	variable T:INTEGER RANGE 1 TO 50000;
	BEGIN
		IF RISING_EDGE(CLK) THEN
			T:=T+1;
			IF T=50000 THEN--50000000
				clk_1k<='1';
				T:=1;
				ELSIF 0<T AND T<25001 THEN--25000001
					clk_1k<='0';
					ELSE
						clk_1k<='1';
			END IF;
		END IF;
	END PROCESS;
	PROCESS(CLK)
	variable T1:INTEGER RANGE 1 TO 50000;
	BEGIN
		IF RISING_EDGE(CLK) THEN
			T1:=T1+1;
			IF T1=50000 THEN--50000000
				clk_100hz<='1';
				T1:=1;
				ELSIF 0<T1 AND T1<25001 THEN--25000001
					clk_100hz<='0';
					ELSE
						clk_100hz<='1';
			END IF;
		END IF;
	END PROCESS;
END BEHAV;