module oled_drive(
	input clk,			//ʱ���ź� 50MHz
	input rst_n,		//������λ
	input ram_rst,		//ram��λ �ߵ�ƽ��λ
	
	input [2:0] count,       //input count_number
	input inputing,             //key_lock
	input input_finish,
	input [2:0] key_num,
	input success,
	
	output oled_rst,	//oled res ��λ�ź�
	output oled_dc,	//oled dc 0��д���� 1��д����
	output oled_sclk,	//oled do ʱ���ź�
	output oled_mosi	//oled d1 �����ź�
);
 
wire clk_1m;			//��Ƶ���1Mʱ��
wire ena_write;		//spiдʹ���ź�
wire [7:0] data;		//spiд������
 
wire init_done;		//��ʼ������ź�
wire [7:0] init_data;//��ʼ�������spi������
wire init_ena_wr;		//��ʼ����spiдʹ���ź�
wire init_oled_dc;
 
wire [7:0] ram_data;	//������ram����
wire [7:0] show_data;//�����spiд������
wire rden;				//ram�Ķ�ʹ���ź�
wire [9:0] rdaddress;//ram����ַ�ź�
wire ram_ena_wr;		//ramʹ��д�ź�
wire ram_oled_dc;		//ramģ���е�oled dc�ź�
 
wire wren;				//ramдʹ���ź�
wire [9:0] wraddress;//ramд��ַ
wire [7:0] wrdata;	//д��ram�е�����
 
//һ���ź�ֻ������һ���ź���������������Ҫѡ��һ��
assign data = init_done ? show_data : init_data;
assign ena_write = init_done ? ram_ena_wr : init_ena_wr;
assign oled_dc = init_done ? ram_oled_dc : init_oled_dc;
 
//ʱ�ӷ�Ƶģ�� ����1M��ʱ��
clk_fenpin clk_fenpin_inst(
	.clk(clk),
	.rst_n(rst_n),
	.clk_1m(clk_1m)
);
 
//spi����ģ��
spi_writebyte spi_writebyte_inst(
	.clk(clk_1m),
	.rst_n(rst_n),
	.ena_write(ena_write),
	.data(data),
	.sclk(oled_sclk),
	.mosi(oled_mosi),
	.write_done(write_done)
);
 
//oled��ʼ��ģ�� ������ʼ������
oled_init oled_init_inst(
	.clk(clk_1m),
	.rst_n(rst_n),
	.write_done(write_done),
	.oled_rst(oled_rst),
	.oled_dc(init_oled_dc),
	.data(init_data),
	.ena_write(init_ena_wr),
	.init_done(init_done)
);
 
//ram��ģ��
ram_read ram_read_inst(
	.clk(clk_1m),
	.rst_n(rst_n),
	.write_done(write_done),
	.init_done(init_done),
	.ram_data(ram_data),
	.rden(rden),
	.rdaddress(rdaddress),
	.ena_write(ram_ena_wr),
	.oled_dc(ram_oled_dc),
	.data(show_data)
);
 
//ramдģ��
ram_write ram_write_inst(
	.clk(clk_1m),
	.rst_n(rst_n),
	.en_ram_wr(1'b1),
	.wren(wren),
	.wraddress(wraddress),
	.data(wrdata),
	.count(count),
	.success(success),
	.inputing(inputing),
	.key_num(key_num),
	.finish_flag(input_finish),
);

//ram ip��
ram_show ram_show_inst(
	.clock(clk_1m),
	.aclr(!ram_rst),
	.data(wrdata),
	.rdaddress(rdaddress),
	.rden(rden),
	.wraddress(wraddress),
	.wren(wren),
	.q(ram_data)
);
endmodule